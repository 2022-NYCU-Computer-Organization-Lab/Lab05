`timescale 1ns/1ps
module Pipeline_CPU(
    clk_i,
    rst_i
);

//I/O port
input         clk_i;
input         rst_i;

// Again, these are the signals TAs forgot to gave us
wire [32-1:0] Imm_4 = 4;
wire [32-1:0] instr;

//Internal Signals
wire [31:0] PC_i;
wire [31:0] PC_o;
wire [31:0] MUXMemtoReg_o;
wire [31:0] ALUResult;
wire [31:0] MUXALUSrc_o;
wire [31:0] Decoder_o;
wire [31:0] RSdata_o;
wire [31:0] RTdata_o;
wire [31:0] Imm_Gen_o;
wire [31:0] ALUSrc1_o;
wire [31:0] ALUSrc2_o;
wire [7:0]  MUX_control_o;

wire [31:0] PC_Add_Immediate;
wire [1:0] ALUOp;
wire PC_write;
wire ALUSrc;
wire RegWrite;
wire Branch;
wire MUXControl; // generated by hazard detection unit
wire Jump;
wire [31:0] SL1_o;
wire [3:0] ALU_Ctrl_o;
wire ALU_zero;
wire Branch_zero;
wire MUXPCSrc;
wire [31:0] DM_o;
wire MemtoReg, MemRead, MemWrite;
wire [1:0] ForwardA;
wire [1:0] ForwardB;
wire [31:0] PC_Add4;

//Pipeline Register Signals
//IFID
wire [31:0] IFID_PC_o;
wire [31:0] IFID_Instr_o;
wire IFID_Write;
wire IFID_Flush;
wire [31:0]IFID_PC_Add4_o;

//IDEXE
wire [31:0] IDEXE_Instr_o;
wire [2:0] IDEXE_WB_o;
wire [1:0] IDEXE_Mem_o;
wire [2:0] IDEXE_Exe_o;
wire [31:0] IDEXE_PC_o;
wire [31:0] IDEXE_RSdata_o;
wire [31:0] IDEXE_RTdata_o;
wire [31:0] IDEXE_ImmGen_o;
wire [3:0] IDEXE_Instr_30_14_12_o;
wire [4:0] IDEXE_Instr_11_7_o;
wire [31:0]IDEXE_PC_add4_o;

//EXEMEM
wire [31:0] EXEMEM_Instr_o;
wire [2:0] EXEMEM_WB_o;
wire [1:0] EXEMEM_Mem_o;
wire [31:0] EXEMEM_PCsum_o;
wire EXEMEM_Zero_o;
wire [31:0] EXEMEM_ALUResult_o;
wire [31:0] EXEMEM_RTdata_o;
wire [4:0]  EXEMEM_Instr_11_7_o;
wire [31:0] EXEMEM_PC_Add4_o;

//MEMWB
wire [2:0] MEMWB_WB_o;
wire [31:0] MEMWB_DM_o;
wire [31:0] MEMWB_ALUresult_o;
wire [4:0]  MEMWB_Instr_11_7_o;
wire [31:0] MEMWB_PC_Add4_o;

assign MUXPCSrc = (Branch & Branch_zero) | Jump;

// IF
MUX_2to1 MUX_PCSrc(
    .data0_i(PC_Add4),
    .data1_i(PC_Add_Immediate),
    .select_i(MUXPCSrc),
    .data_o(pc_i)
);

ProgramCounter PC(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .pc_i(pc_i),
    .pc_o(pc_o)
);

Adder PC_plus_4_Adder(
    .src1_i(pc_o),
    .src2_i(Imm_4),
    .sum_o(PC_Add4)
);

Instr_Memory IM(
    .addr_i(pc_o),
    instr_o(instr)
);

IFID_register IFtoID(
);

// ID
Hazard_detection Hazard_detection_obj(
);

MUX_2to1 MUX_control(
);

Decoder Decoder(
);

Reg_File RF(
);

Imm_Gen ImmGen(
);

Shift_Left_1 SL1(
);

Adder Branch_Adder(
);

IDEXE_register IDtoEXE(
);

// EXE
MUX_2to1 MUX_ALUSrc(
);

ForwardingUnit FWUnit(
);

MUX_3to1 MUX_ALU_src1(
);

MUX_3to1 MUX_ALU_src2(
);

ALU_Ctrl ALU_Ctrl(
);

alu alu(
);

EXEMEM_register EXEtoMEM(
);

// MEM
Data_Memory Data_Memory(
);

MEMWB_register MEMtoWB(
);

// WB
MUX_3to1 MUX_MemtoReg(
);

endmodule
